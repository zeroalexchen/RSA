module moutmul(x,y,z)
    input   [2047,0] x;
    input   [2047,0] y;
    reg     [2047,0] i;
    reg     [2047,0] temp1;
    output  [2047,0] z;

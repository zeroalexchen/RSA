module MONT_REDC(t,result);
	input [2047:0] t;
	
	output reg [2047:0] result;


endmodule
`timescale 1ns/1ns
`include "RSA_TOP.V"
module exp_top;
	reg 	[2047:0] 	c;
	reg  	[2047:0] 	e;
	reg 	[2047:0] 	n;
	reg 				enable;
	reg					clk;
	reg					sys_rst;

	wire	 [2047:0]	result;
	wire 				finish;

	RSA_TOP rsa_top_u(.c(c),.e(e),.n(n),.enable(enable),.clk(clk),.sys_rst(sys_rst),.result(result),.finish(finish));

initial begin
	$dumpfile("test.vcd");
	$dumpvars(0,rsa_top_u);
/*	c = 'h3DB5F1F063E96712232D9F5464294F0CD1F19AD562B45627C8EBEBAB9FF8D416F06A74BDFF06036227B78CC421A6FF0241D34447174C6290FDBF608302FD6780B43B76E906890256CDAF6A0986260E3419B5970A8EBD70A0C71CC25E6BA6E85E3DD22513225B334C20D9FCA9325F337C23769E7FB9A0EE9138FE6BD53888082AB35F5A30F7B1F08F4549D284A0D905528723140A803680C47DE8179C8E914E23B08FB5762D4792EDF64BE02B9B85C7E9F68BCE154E52D5620E5877D3DF567B686AC88E08B5D9DF0D4E6C67E0F692C30AC2794285B2FDB92DB21ECF0F98354640F89E1C8E83CE2B684B58B4B9F72C1F5B7EE6BEEAD13510EF8A95E8690B8B76E7;
	e = 'h37BA4B62B92169699F52DDDCCD81C0B4E2D216B3328A45B93D8DD9E7B9EFCB02B7C2C50D7195C6BBB9877F4C32F1C002178774377E234F8B4CD7FE62F94EF47D4CA47ADA70ECDDB6A1370A6D6D1ACBA0DFB0DB3F6B2EC334AC92F0FB492C10E7E6E5EEABCA5196C9ACCB55B6DCDCF07DEEFFB2DCFEBA70E8D405EB9DCB3A8A7DCB570D84C13723DB389740922BA681343FE8605775062B090270B6CB7BF0C2BF8096FBC27E665183B1DE78F6EF3A66B83E656326472F28201A7ACB4FE3224F9E01AEAC93A9E5D60F4977B572D75F109DE5056AB4FC8B4D4BD884E09AFE8B9D844B2969D7E7878AAC595ADF411B7DE2F2FC147751B3D15DBA7D83B0C1E96729FE;
	e = 'hf;
	n = 'hDE68957574712E6D38EFAAA4C06E769AD854B1F70686AD11DFB7DADAA6E97B43AB78B6C1F650B578FB3F0ECB99AC32A3758FD99782DEDCE8C4874ED2F2120933C46B1D3DD71B0F0229BB6994397AD11B5F1A329E02A0DC18DED4E34D611855EFAAEBB0CF83D82B50EEFE032D6FD6CFE071FE9CDACFFCE74F115503087BAE630DD7369DB06A484F7319D61DC0D93E0D2B090563C93F4D17DB4165B93E1B9D967167849D330DB415572F69E79AFB47B8860137E0AB30ED169583F2FE5DE170795FEDB22C69368D6FB3D2FCC8D0E7AD1A3458174B8498A0925DA44AFDC16510DBC40158A8545FE43CA8F0ED066BB16477DEABBD3BABF8398ECC2D45483E37865071;*/

	c = 'h161018d2ec6c64b175726b05844a5973cbffbde17ad56ddbdeed1decc249cfed4773033bf3eee49b0b287aed4e63cf04e04008e1470751a9f8618050c6d5185e8b0bd7260deedca880aaaac19622dccfb8a525826294d4e58eb4219c5046f9d56ea39541eaf35ffa5e86d657b0cc70a6f487453fd8a3c47972540eb2b7bc4b9473333cdb94e3d64baf682ed501d809bee3bc6490745bd32dac402e7a0ab811220a1f03d10a81911a38e1f5ee1d31bb97f5706e5608bf0850df9c2766373f9e838bbd7c41c8ee0b1151a4ff15f8892072dfe4d94fce635e11f750121f0d32ac5206ea2d3b2297dfe35d416cec1a5d4187edc58456452ed0a021aa2123d0b83c87;
	e = 'h2474fe4fb0268a6f2efd9ed7541abde46cbb54e7dbbf16469ec41254266b0e70e6182ba87d07cc039d275fd463f9bf6bb4f311a3c4f72f413a6a768101618dc15454c6df889897b16a402ef1cbcfa23c1bcfca525d2dc49bed3eb268f7579d53e4fa6a7e8db78809ebeb1e4120d60d92b6ae30f821f3f65fb0af5b28b39658b32cbaad6d66da6f325849fcab656d4ddb8a382701d5e15cbd35faa9fa388c91724e696be3d76b4462cd61388e7cc756c8e1d025f79eaa438301ba6363544c80a127a3d79c3c6a0309ae649f55b30c8c4a9a9e358335ec6e2bc01e94938cb1c50bd8aaa30a1238b9c7c1c988f96c8d447a250aa025c493a865bc7169d97d06af71;
	n = 'h81c82370cec71b5cb6bab156013264b841a168eb66b0f6269db9c3c3b758c1bb0946a2ed03c229b550e3572f230b330da90bbe928b5fc1991127b2f4ca63626851f5dda144b900aae5cbe61b9238dfc374c6e0cc591bb26015baa2778e511b2a1c2d44d87bc9ae88b7d850eef07139627b700ba844eabaaa592fa46833c930502c2a09ca601dc5f28821465063643abc67d8df06a84df9805f2eeba760ba7e3e8f3b77ae4f6d0e223c30942228b304c636fbaad770080fa9ebb21a088b0ff370f9dd5b0342a9d44e5183c28ddb0d36aff49a2577a5f1776a66db45247ab309b7879c6fe9c30765d67087111c353c23ef77dc7902d931ec5bef39a8dcf0891a93;

/*
	c = 59855131;
	e = 787;
	n = 5959137;
*/
	enable = 1;
	sys_rst = 1;
	#5;
	sys_rst = 0;
	#5;
	wait(finish)
	#50;
		$display("result = %d\nfinish = %b",result,finish);
		$display("time = %d ns",$realtime);
	$finish;

end

always begin
	clk = 0;
	#5;
	clk = 1;
	#5;
end

endmodule